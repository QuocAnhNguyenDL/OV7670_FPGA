module CAM_SDRAM_VGA
(
	input CLOCK_50,
	
	//-------------CAM_SIGNALS------------------
	output				CMOS_SCLK,		//cmos i2c clock
	inout					CMOS_SDAT,		//cmos i2c data
	input					CMOS_VSYNC,		//cmos vsync
	input					CMOS_HREF,		//cmos hsync refrence
	input					CMOS_PCLK,		//cmos pxiel clock
	output				CMOS_XCLK,		//cmos externl clock
	input		[7 :0]	CMOS_DB,		//cmos data
	
	//-----------SDRAM CONTROLLER SIGNALS--------
	output				S_CLK,		//sdram clock
	output				S_CKE,		//sdram clock enable
	output				S_NCS,		//sdram chip select
	output				S_NWE,		//sdram write enable
	output				S_NCAS,	//sdram column address strobe
	output				S_NRAS,	//sdram row address strobe
	output	[1 :0] 	S_DQM,		//sdram data enable 
	output	[1 :0]	S_BA,		//sdram bank address
	output	[11:0]	S_A,		//sdram address
	inout		[15:0]	S_DB,		//sdram data
	
	//------------VGA SIGNALS----------			
	output			VGA_HS,			//horizontal sync 
	output			VGA_VS,			//vertical sync
	output 			VGA_BLANK,
	output	[15:0]VGAD,		//VGA data
	output         VGA_CLK
);


//-------------CONTROL--------------
wire	clk_vga;		
wire	clk_ref;		
wire	clk_refout;		
wire	sys_rst_n;		
system_ctrl	my_system_ctrl
(
	.clk					(CLOCK_50	),			
	.rst_n				(rst_n		),		
	
	.sys_rst_n			(sys_rst_n	),	
	.clk_c0				(clk_vga		),		
	.clk_c1				(clk_ref		),		
	.clk_c2				(clk_refout	)	
);
assign VGA_CLK = clk_vga;
assign rst_n = 1'b1;

//------------CAM OV7670------------
wire 			sys_we;
wire [15:0] sys_data_in;
wire 			frame_valid;
CAM cam
(
	.clk_vga				(clk_vga		),
	.sys_rst_n			(sys_rst_n	),
	
	.sdram_init_done	(sdram_init_done),
	
	.CMOS_SCLK			(CMOS_SCLK	),		//cmos i2c clock
	.CMOS_SDAT			(CMOS_SDAT	),		//cmos i2c data
	.CMOS_VSYNC			(CMOS_VSYNC	),		//cmos vsync
	.CMOS_HREF			(CMOS_HREF	),		//cmos hsync refrence
	.CMOS_PCLK			(CMOS_PCLK	),		//cmos pxiel clock
	.CMOS_XCLK			(CMOS_XCLK	),		//cmos externl clock
	.CMOS_DB				(CMOS_DB		),		//cmos data
	
	.CMOS_oCLK			(sys_we		),
	.CMOS_oDATA			(sys_data_in),
	.CMOS_VALID			(frame_valid)
);

//----------------SDRAM CONTROLLER----------------
wire sdram_init_done;
wire sys_rd;
wire [15:0] sys_data_out;
wire vga_frame;
SDRAM_TOP SDRAM
(
	//global clock
	.clk_vga				(clk_vga),		//vga clock
	.clk_ref				(clk_ref),		//sdram ctrl clock
	.clk_refout			(clk_refout),		//sdram clock output
	.rst_n				(rst_n),			//global reset

	//sdram control
	.sdram_clk			(S_CLK),		//sdram clock
	.sdram_cke			(S_CKE),		//sdram clock enable
	.sdram_cs_n			(S_NCS),		//sdram chip select
	.sdram_we_n			(S_NWE),		//sdram write enable
	.sdram_cas_n		(S_NCAS),		//sdram column address strobe
	.sdram_ras_n		(S_NRAS),		//sdram row address strobe
	.sdram_udqm			(S_DQM[1]),		//sdram data enable (H:8)
	.sdram_ldqm			(S_DQM[0]),		//sdram data enable (L:8)
	.sdram_ba			(S_BA),			//sdram bank address
	.sdram_addr			(S_A),		//sdram address
	.sdram_data			(S_DB),		//sdram data
		
	//user interface read
	.clk_write			(clk_vga),		//fifo write clock
	.sys_we				(sys_we),			//fifo write enable
	.sys_data_in		(sys_data_in),	//fifo data input
	.sdram_init_done	(sdram_init_done),//sdram init done
	.frame_valid		(frame_valid),		//frame valid
	
	//user interface write
	.sys_rd				(sys_rd),        		//fifo read enable
	.sys_data_out		(sys_data_out),  		//fifo data output
	.vga_framesync		(vga_framesyn)		//vga frame sync
);

VGA vga
(  	
	//global clock
	.clk					(clk_vga),			
	.rst_n				(rst_n),     		
	
	//vga interface
	.vga_blank			(VGA_BLANK),				
	.vga_hs				(VGA_HS),	    	
	.vga_vs				(VGA_VS),	    				
	.vga_rgb				(VGAD),		
	
	//user interface
	.vga_request(sys_rd),	//vga data request
	.vga_framesync	(vga_framesyn),	//vga frame sync
	.vga_data(sys_data_out)		//vga data
);	 

endmodule